`include "FullAdder_GL.v"

module complexrhs_port_test_pass (
    input wire [1:0] in0,
    input wire [1:0] in1,
    input wire cin,
    output wire [1:0] sum,
    output wire cout
);

    

endmodule

