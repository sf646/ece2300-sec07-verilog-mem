
module primonly_test_pass(
    input logic a,
    input logic b,
    output logic y
);

assign y = a & b;

endmodule

