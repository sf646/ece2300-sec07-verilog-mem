
module nospblk_test_pass(
    input logic a,
    input logic b,
    output logic y
);

and(y, a, b);

endmodule

