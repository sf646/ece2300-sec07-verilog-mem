//========================================================================
// RegfileStruct1r1w_4x4b_RTL-test
//========================================================================

`include "ece2300/ece2300-test.v"

// ece2300-lint
`include "mem/RegfileStruct1r1w_4x4b_RTL.v"

module Top();

  //----------------------------------------------------------------------
  // Setup
  //----------------------------------------------------------------------

  logic clk;
  logic rst;

  TestUtilsClkRst t( .* );

  `ECE2300_UNUSED( rst );

  //----------------------------------------------------------------------
  // Instantiate design under test
  //----------------------------------------------------------------------

  logic       wen;
  logic [1:0] waddr;
  logic [3:0] wdata;
  logic [1:0] raddr;
  logic [3:0] rdata;

  RegfileStruct1r1w_4x4b_RTL dut ( .* );

  //----------------------------------------------------------------------
  // Include test cases
  //----------------------------------------------------------------------

  `include "mem/test/Regfile1r1w_4x4b-test-cases.v"

endmodule

