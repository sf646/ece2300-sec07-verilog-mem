
module complexlhs_test_pass(
    input logic a,
    input logic b,
    output logic y,
    output logic v
);

assign y = a;
assign v = b;

endmodule

